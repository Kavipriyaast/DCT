// Module: clock_gating
// Description: This module implements a simple clock gating mechanism. 
//              Clock gating is a technique used to reduce power consumption 
//              by disabling the clock signal to certain parts of a circuit 
//              when they are not in use. This is achieved by ANDing the 
//              clock signal with an enable signal.

module clock_gating (
    input clk,        // Input clock signal
    input enable,     // Enable signal to control clock gating
    output gated_clk  // Output gated clock signal
);

    // The gated clock is generated by ANDing the input clock with the enable signal.
    // When 'enable' is high, 'gated_clk' follows 'clk'.
    // When 'enable' is low, 'gated_clk' is held low, effectively disabling the clock.
    assign gated_clk = clk & enable;

endmodule
